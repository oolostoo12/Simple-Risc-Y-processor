`timescale 1ns/ 100ps
package phasepackage;
   typedef enum [1:0] {FETCH,DECODE,EXECUTE,UPDATE}STATE;
endpackage // phasepackage
   